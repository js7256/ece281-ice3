(Shearer, Joseph R C4C USAF USAFA CW/CS28             ( S h e a r e r ,   J o s e p h   R   C 4 C   U S A F   U S A F A   C W / C S 2 8           -ˤ    J= ��T